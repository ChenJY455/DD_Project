module top(

    );
    
endmodule